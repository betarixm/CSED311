`include "env.v"

module dmac(clk, reset_n);
    input clk;
    input reset_n;
endmodule